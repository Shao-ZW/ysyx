module ALU(

);


endmodule