module Control(

);


endmodule